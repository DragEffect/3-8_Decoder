interface add_if(input logic clk, reset);
  logic [2:0] ip;
  logic [7:0] out;
  
endinterface
